.SUBCKT modulator 1 2 3
E1 4 0 2 0 0.5
V1 5 0 dc=-0.5V
B1 3 0 V=v(4,5)*v(1)
.ENDS